
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41.500.3.38
#
# TECH LIB NAME: tsmc18
# TECH FILE NAME: techfile.cds
#******

VERSION 5.4 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "|" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 100  ;
END UNITS

MACRO FIR_Fliter
    CLASS CORE ;
    FOREIGN FIR_Fliter 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 120.13 BY 120.13 ;
    SYMMETRY X Y ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 118 0.2 118.2 ;
        END
        AntennaGateArea 0.0 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 113 0.2 113.2 ;
        END
        AntennaGateArea 0.0 ;
    END SE
    PIN A[0]
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 108 0.2 108.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[0]
    PIN Signal_Noise[1]
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 103 0.2 103.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[1]
    PIN Signal_Noise[2]
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 98 0.2 98.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[2]
    PIN Signal_Noise[3]
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 93 0.2 93.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[3]
    PIN Signal_Noise[4]
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 88 0.2 88.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[4]
    PIN Signal_Noise[5]
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 83 0.2 83.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[5]
    PIN Signal_Noise[6]
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 78 0.2 78.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[6]
    PIN Signal_Noise[7]
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 73 0.2 73.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[7]
   
 PIN Signal_Noise[8]
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 43 0.2 43.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[8]
    PIN Signal_Noise[9]
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 38 0.2 38.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[9]
    PIN Signal_Noise[10]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 33 0.2 33.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[10]
    PIN Signal_Noise[11]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 28 0.2 28.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[11]
    PIN Signal_Noise[12]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 23 0.2 23.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[12]
    PIN Signal_Noise[13]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 18 0.2 18.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[13]
    PIN Signal_Noise[14]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 13 0.2 13.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[14]
    PIN Signal_Noise[15]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 8 0.2 8.2 ;
        END
        AntennaGateArea 0.0 ;
    END Signal_Noise[15] 
   PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 68 0.2 68.2 ;
        END
        AntennaGateArea 0.0 ;
    END CLK
    PIN scan_clk
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 58 0.2 58.2 ;
        END
        AntennaGateArea 0.0 ;
    END scan_clk
    PIN scan_rst
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 53 0.2 53.2 ;
        END
        AntennaGateArea 0.0 ;
    END scan_rst
    PIN test_mode
        DIRECTION INPUT ;
        PORT
        LAYER METAL3 ;
        RECT  0.00 48 0.2 48.2 ;
        END
        AntennaGateArea 0.0 ;
    END test_mode
  
    PIN Fliter_Signal[0]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL5 ;
        RECT  25 0.0 25.2 0.2 ;
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[0]
    PIN Fliter_Signal[1]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL5 ;
        RECT  30 0.0 30.2 0.2 ;
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[1]
    PIN Fliter_Signal[2]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL5 ;
        RECT  35 0.0 35.2 0.2 ;
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[2]
    PIN Fliter_Signal[3]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL5 ;
        RECT  40 0.0 40.2 0.2 ;
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[3]
    PIN Fliter_Signal[4]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL5 ;
        RECT  45 0.0 45.2 0.2 ;
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[4]
    PIN Fliter_Signal[5]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL5 ;
        RECT  50 0.0 50.2 0.2 ;
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[5]
    PIN Fliter_Signal[6]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL5 ;
        RECT  55 0.0 55.2 0.2 ;
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[6]
    PIN Fliter_Signal[7]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL5 ;
        RECT  60 0.0 60.2 0.2 ;
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[7]
    PIN Fliter_Signal[8]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL3 ;
        RECT  119.83 108 120.13 108.2 ; 
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[8]
    PIN Fliter_Signal[9]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL3 ;
        RECT  119.83 103 120.13 103.2 ; 
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[9]
    PIN Fliter_Signal[10]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL3 ;
        RECT  119.83 98 120.13 98.2 ; 
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[10]
    PIN Fliter_Signal[11]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL3 ;
        RECT  119.83 93 120.13 93.2 ; 
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[11]
    PIN Fliter_Signal[12]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL3 ;
        RECT  119.83 88 120.13 88.2 ; 
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[12]
    PIN Fliter_Signal[13]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL3 ;
        RECT  119.83 83 120.13 83.2 ; 
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[13]
    PIN Fliter_Signal[14]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL3 ;
        RECT  119.83 78 120.13 78.2 ; 
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[14]
    PIN Fliter_Signal[15]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL3 ;
        RECT  119.83 73 120.13 73.2 ; 
        END
        AntennaDiffArea 0.575 ;
    END Fliter_Signal[15]
    PIN SO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL3 ;
        RECT  70 0.0 70.2 0.2 ;
        END
        AntennaDiffArea 0.575 ;
    END SO
END FIR_Fliter

END LIBRARY

